* C:\Users\zelle\Desktop\���\2����\3���\�����\����7\Lab7.sch

* Schematics Version 9.2
* Mon Dec 11 21:35:27 2023



** Analysis setup **
.tran 20ns 50us


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Lab7.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
